goodhands
R1_M 12 14 1000
CRing 9 18 1µF IC=0
R1_M 12 9 1000
R1_M 12 16 1000
R7 2 0 220
R8 3 0 220
R5 4 0 220
R1_M 12 15 1000
R6 1 0 220

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
